`timescale 1ns/1ns

module tb_avoid_latch()
{
    reg in1,in2,in3;
    wire [7:0]out
};

initial  begin
       

end
    

    avoid_latch avoid_latch_inst
    (
        .in1(in1),
        .in2(in2),
        .in3(in3),
        .out(out)

    );

end